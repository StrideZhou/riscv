`include "mem.vh"
module dmem_mod (
	input        clk,
	input		 nrst,
	input		 stall,
	input [31:0] inst
	
//todo: depands on alu_mod
);



endmodule